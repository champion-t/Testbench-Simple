package my_pkg;
    `include "packet.sv"
    `include "driver.sv"
    `include "monitor.sv"
    `include "scoreboard.sv"
    `include "environment.sv"
    `include "test.sv"
endpackage